  LIBRARY ieee; USE ieee.std_logic_1164.ALL; LIBRARY XilinxCoreLib; ENTITY MAC01_2_75F243352369479695E2AED5F4206BF1 IS   PORT (     clk : in std_logic := '0';     ce : IN STD_LOGIC;     sclr : IN STD_LOGIC;     bypass : IN STD_LOGIC;     a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     s : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)   ); END MAC01_2_75F243352369479695E2AED5F4206BF1;  ARCHITECTURE MAC01_2_75F243352369479695E2AED5F4206BF1_a OF MAC01_2_75F243352369479695E2AED5F4206BF1 IS COMPONENT wrapped_MAC01_2_75F243352369479695E2AED5F4206BF1   PORT (     clk : IN STD_LOGIC;     ce : IN STD_LOGIC;     sclr : IN STD_LOGIC;     bypass : IN STD_LOGIC;     a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     s : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)   ); END COMPONENT;    FOR ALL : wrapped_MAC01_2_75F243352369479695E2AED5F4206BF1 USE ENTITY XilinxCoreLib.xbip_multaccum_v2_0(behavioral)     GENERIC MAP (       c_a_type => 0,       c_a_width => 32,       c_accum_mode => 0,       c_accum_width => 64,       c_b_type => 0,       c_b_width => 32,       c_bypass_low => 0,       c_ce_overrides_sclr => 0,       c_has_bypass => 1,       c_latency => -1,       c_out_width => 36,       c_round_type => 0,       c_use_dsp48 => 1,       c_verbosity => 0,       c_xdevicefamily => "spartan6"     ); BEGIN U0 : wrapped_MAC01_2_75F243352369479695E2AED5F4206BF1   PORT MAP (     clk => clk,     ce => ce,     sclr => sclr,     bypass => bypass,     a => a,     b => b,     s => s   );  END MAC01_2_75F243352369479695E2AED5F4206BF1_a; 
configuration conf_75F243352369479695E2AED5F4206BF1 of MAC01_2_75F243352369479695E2AED5F4206BF1 is
  for MAC01_2_75F243352369479695E2AED5F4206BF1_a end for; 
end conf_75F243352369479695E2AED5F4206BF1; 